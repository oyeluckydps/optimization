// Float_4E3M Adder - Behavioral Verilog
// Generated from truth table

module float_4e3m_adder(
    input [15:0] operands,  // {op1[7:0], op2[7:0]}
    output reg [7:0] result
);

always @(*) begin
    case (operands)
        16'b0000000000000000: result = 8'b00000111;
        16'b0000000000000001: result = 8'b00000111;
        16'b0000000000000010: result = 8'b00000111;
        16'b0000000000000011: result = 8'b00000111;
        16'b0000000000000100: result = 8'b00000111;
        16'b0000000000000101: result = 8'b00000111;
        16'b0000000000000110: result = 8'b00000111;
        16'b0000000000000111: result = 8'b00000111;
        16'b0000000000001000: result = 8'b00000100;
        16'b0000000000001001: result = 8'b00000100;
        16'b0000000000001010: result = 8'b00000101;
        16'b0000000000001011: result = 8'b00000101;
        16'b0000000000001100: result = 8'b00000110;
        16'b0000000000001101: result = 8'b00000110;
        16'b0000000000001110: result = 8'b00000111;
        16'b0000000000001111: result = 8'b00000111;
        16'b0000000100000000: result = 8'b00000111;
        16'b0000000100000001: result = 8'b00000111;
        16'b0000000100000010: result = 8'b00000111;
        16'b0000000100000011: result = 8'b00000111;
        16'b0000000100000100: result = 8'b00000111;
        16'b0000000100000101: result = 8'b00000111;
        16'b0000000100000110: result = 8'b00000111;
        16'b0000000100000111: result = 8'b00000111;
        16'b0000000100001000: result = 8'b00000101;
        16'b0000000100001001: result = 8'b00000101;
        16'b0000000100001010: result = 8'b00000110;
        16'b0000000100001011: result = 8'b00000110;
        16'b0000000100001100: result = 8'b00000111;
        16'b0000000100001101: result = 8'b00000111;
        16'b0000000100001110: result = 8'b00000111;
        16'b0000000100001111: result = 8'b00000111;
        16'b0000001000000000: result = 8'b00000111;
        16'b0000001000000001: result = 8'b00000111;
        16'b0000001000000010: result = 8'b00000111;
        16'b0000001000000011: result = 8'b00000111;
        16'b0000001000000100: result = 8'b00000111;
        16'b0000001000000101: result = 8'b00000111;
        16'b0000001000000110: result = 8'b00000111;
        16'b0000001000000111: result = 8'b00000111;
        16'b0000001000001000: result = 8'b00000110;
        16'b0000001000001001: result = 8'b00000110;
        16'b0000001000001010: result = 8'b00000111;
        16'b0000001000001011: result = 8'b00000111;
        16'b0000001000001100: result = 8'b00000111;
        16'b0000001000001101: result = 8'b00000111;
        16'b0000001000001110: result = 8'b00000111;
        16'b0000001000001111: result = 8'b00000111;
        16'b0000001100000000: result = 8'b00000111;
        16'b0000001100000001: result = 8'b00000111;
        16'b0000001100000010: result = 8'b00000111;
        16'b0000001100000011: result = 8'b00000111;
        16'b0000001100000100: result = 8'b00000111;
        16'b0000001100000101: result = 8'b00000111;
        16'b0000001100000110: result = 8'b00000111;
        16'b0000001100000111: result = 8'b00000111;
        16'b0000001100001000: result = 8'b00000111;
        16'b0000001100001001: result = 8'b00000111;
        16'b0000001100001010: result = 8'b00000111;
        16'b0000001100001011: result = 8'b00000111;
        16'b0000001100001100: result = 8'b00000111;
        16'b0000001100001101: result = 8'b00000111;
        16'b0000001100001110: result = 8'b00000111;
        16'b0000001100001111: result = 8'b00000111;
        16'b0000010000000000: result = 8'b00000111;
        16'b0000010000000001: result = 8'b00000111;
        16'b0000010000000010: result = 8'b00000111;
        16'b0000010000000011: result = 8'b00000111;
        16'b0000010000000100: result = 8'b00000111;
        16'b0000010000000101: result = 8'b00000111;
        16'b0000010000000110: result = 8'b00000111;
        16'b0000010000000111: result = 8'b00000111;
        16'b0000010000001000: result = 8'b00000111;
        16'b0000010000001001: result = 8'b00000111;
        16'b0000010000001010: result = 8'b00000111;
        16'b0000010000001011: result = 8'b00000111;
        16'b0000010000001100: result = 8'b00000111;
        16'b0000010000001101: result = 8'b00000111;
        16'b0000010000001110: result = 8'b00000111;
        16'b0000010000001111: result = 8'b00000111;
        16'b0000010100000000: result = 8'b00000111;
        16'b0000010100000001: result = 8'b00000111;
        16'b0000010100000010: result = 8'b00000111;
        16'b0000010100000011: result = 8'b00000111;
        16'b0000010100000100: result = 8'b00000111;
        16'b0000010100000101: result = 8'b00000111;
        16'b0000010100000110: result = 8'b00000111;
        16'b0000010100000111: result = 8'b00000111;
        16'b0000010100001000: result = 8'b00000111;
        16'b0000010100001001: result = 8'b00000111;
        16'b0000010100001010: result = 8'b00000111;
        16'b0000010100001011: result = 8'b00000111;
        16'b0000010100001100: result = 8'b00000111;
        16'b0000010100001101: result = 8'b00000111;
        16'b0000010100001110: result = 8'b00000111;
        16'b0000010100001111: result = 8'b00000111;
        16'b0000011000000000: result = 8'b00000111;
        16'b0000011000000001: result = 8'b00000111;
        16'b0000011000000010: result = 8'b00000111;
        16'b0000011000000011: result = 8'b00000111;
        16'b0000011000000100: result = 8'b00000111;
        16'b0000011000000101: result = 8'b00000111;
        16'b0000011000000110: result = 8'b00000111;
        16'b0000011000000111: result = 8'b00000111;
        16'b0000011000001000: result = 8'b00000111;
        16'b0000011000001001: result = 8'b00000111;
        16'b0000011000001010: result = 8'b00000111;
        16'b0000011000001011: result = 8'b00000111;
        16'b0000011000001100: result = 8'b00000111;
        16'b0000011000001101: result = 8'b00000111;
        16'b0000011000001110: result = 8'b00000111;
        16'b0000011000001111: result = 8'b00000111;
        16'b0000011100000000: result = 8'b00000111;
        16'b0000011100000001: result = 8'b00000111;
        16'b0000011100000010: result = 8'b00000111;
        16'b0000011100000011: result = 8'b00000111;
        16'b0000011100000100: result = 8'b00000111;
        16'b0000011100000101: result = 8'b00000111;
        16'b0000011100000110: result = 8'b00000111;
        16'b0000011100000111: result = 8'b00000111;
        16'b0000011100001000: result = 8'b00000111;
        16'b0000011100001001: result = 8'b00000111;
        16'b0000011100001010: result = 8'b00000111;
        16'b0000011100001011: result = 8'b00000111;
        16'b0000011100001100: result = 8'b00000111;
        16'b0000011100001101: result = 8'b00000111;
        16'b0000011100001110: result = 8'b00000111;
        16'b0000011100001111: result = 8'b00000111;
        16'b0000100000000000: result = 8'b00000100;
        16'b0000100000000001: result = 8'b00000101;
        16'b0000100000000010: result = 8'b00000110;
        16'b0000100000000011: result = 8'b00000111;
        16'b0000100000000100: result = 8'b00000111;
        16'b0000100000000101: result = 8'b00000111;
        16'b0000100000000110: result = 8'b00000111;
        16'b0000100000000111: result = 8'b00000111;
        16'b0000100000001000: result = 8'b00000000;
        16'b0000100000001001: result = 8'b00000000;
        16'b0000100000001010: result = 8'b00000001;
        16'b0000100000001011: result = 8'b00000001;
        16'b0000100000001100: result = 8'b00000010;
        16'b0000100000001101: result = 8'b00000010;
        16'b0000100000001110: result = 8'b00000011;
        16'b0000100000001111: result = 8'b00000011;
        16'b0000100100000000: result = 8'b00000100;
        16'b0000100100000001: result = 8'b00000101;
        16'b0000100100000010: result = 8'b00000110;
        16'b0000100100000011: result = 8'b00000111;
        16'b0000100100000100: result = 8'b00000111;
        16'b0000100100000101: result = 8'b00000111;
        16'b0000100100000110: result = 8'b00000111;
        16'b0000100100000111: result = 8'b00000111;
        16'b0000100100001000: result = 8'b00000000;
        16'b0000100100001001: result = 8'b00000001;
        16'b0000100100001010: result = 8'b00000001;
        16'b0000100100001011: result = 8'b00000010;
        16'b0000100100001100: result = 8'b00000010;
        16'b0000100100001101: result = 8'b00000011;
        16'b0000100100001110: result = 8'b00000011;
        16'b0000100100001111: result = 8'b00000100;
        16'b0000101000000000: result = 8'b00000101;
        16'b0000101000000001: result = 8'b00000110;
        16'b0000101000000010: result = 8'b00000111;
        16'b0000101000000011: result = 8'b00000111;
        16'b0000101000000100: result = 8'b00000111;
        16'b0000101000000101: result = 8'b00000111;
        16'b0000101000000110: result = 8'b00000111;
        16'b0000101000000111: result = 8'b00000111;
        16'b0000101000001000: result = 8'b00000001;
        16'b0000101000001001: result = 8'b00000001;
        16'b0000101000001010: result = 8'b00000010;
        16'b0000101000001011: result = 8'b00000010;
        16'b0000101000001100: result = 8'b00000011;
        16'b0000101000001101: result = 8'b00000011;
        16'b0000101000001110: result = 8'b00000100;
        16'b0000101000001111: result = 8'b00000100;
        16'b0000101100000000: result = 8'b00000101;
        16'b0000101100000001: result = 8'b00000110;
        16'b0000101100000010: result = 8'b00000111;
        16'b0000101100000011: result = 8'b00000111;
        16'b0000101100000100: result = 8'b00000111;
        16'b0000101100000101: result = 8'b00000111;
        16'b0000101100000110: result = 8'b00000111;
        16'b0000101100000111: result = 8'b00000111;
        16'b0000101100001000: result = 8'b00000001;
        16'b0000101100001001: result = 8'b00000010;
        16'b0000101100001010: result = 8'b00000010;
        16'b0000101100001011: result = 8'b00000011;
        16'b0000101100001100: result = 8'b00000011;
        16'b0000101100001101: result = 8'b00000100;
        16'b0000101100001110: result = 8'b00000100;
        16'b0000101100001111: result = 8'b00000101;
        16'b0000110000000000: result = 8'b00000110;
        16'b0000110000000001: result = 8'b00000111;
        16'b0000110000000010: result = 8'b00000111;
        16'b0000110000000011: result = 8'b00000111;
        16'b0000110000000100: result = 8'b00000111;
        16'b0000110000000101: result = 8'b00000111;
        16'b0000110000000110: result = 8'b00000111;
        16'b0000110000000111: result = 8'b00000111;
        16'b0000110000001000: result = 8'b00000010;
        16'b0000110000001001: result = 8'b00000010;
        16'b0000110000001010: result = 8'b00000011;
        16'b0000110000001011: result = 8'b00000011;
        16'b0000110000001100: result = 8'b00000100;
        16'b0000110000001101: result = 8'b00000100;
        16'b0000110000001110: result = 8'b00000101;
        16'b0000110000001111: result = 8'b00000101;
        16'b0000110100000000: result = 8'b00000110;
        16'b0000110100000001: result = 8'b00000111;
        16'b0000110100000010: result = 8'b00000111;
        16'b0000110100000011: result = 8'b00000111;
        16'b0000110100000100: result = 8'b00000111;
        16'b0000110100000101: result = 8'b00000111;
        16'b0000110100000110: result = 8'b00000111;
        16'b0000110100000111: result = 8'b00000111;
        16'b0000110100001000: result = 8'b00000010;
        16'b0000110100001001: result = 8'b00000011;
        16'b0000110100001010: result = 8'b00000011;
        16'b0000110100001011: result = 8'b00000100;
        16'b0000110100001100: result = 8'b00000100;
        16'b0000110100001101: result = 8'b00000101;
        16'b0000110100001110: result = 8'b00000101;
        16'b0000110100001111: result = 8'b00000110;
        16'b0000111000000000: result = 8'b00000111;
        16'b0000111000000001: result = 8'b00000111;
        16'b0000111000000010: result = 8'b00000111;
        16'b0000111000000011: result = 8'b00000111;
        16'b0000111000000100: result = 8'b00000111;
        16'b0000111000000101: result = 8'b00000111;
        16'b0000111000000110: result = 8'b00000111;
        16'b0000111000000111: result = 8'b00000111;
        16'b0000111000001000: result = 8'b00000011;
        16'b0000111000001001: result = 8'b00000011;
        16'b0000111000001010: result = 8'b00000100;
        16'b0000111000001011: result = 8'b00000100;
        16'b0000111000001100: result = 8'b00000101;
        16'b0000111000001101: result = 8'b00000101;
        16'b0000111000001110: result = 8'b00000110;
        16'b0000111000001111: result = 8'b00000110;
        16'b0000111100000000: result = 8'b00000111;
        16'b0000111100000001: result = 8'b00000111;
        16'b0000111100000010: result = 8'b00000111;
        16'b0000111100000011: result = 8'b00000111;
        16'b0000111100000100: result = 8'b00000111;
        16'b0000111100000101: result = 8'b00000111;
        16'b0000111100000110: result = 8'b00000111;
        16'b0000111100000111: result = 8'b00000111;
        16'b0000111100001000: result = 8'b00000011;
        16'b0000111100001001: result = 8'b00000100;
        16'b0000111100001010: result = 8'b00000100;
        16'b0000111100001011: result = 8'b00000101;
        16'b0000111100001100: result = 8'b00000101;
        16'b0000111100001101: result = 8'b00000110;
        16'b0000111100001110: result = 8'b00000110;
        16'b0000111100001111: result = 8'b00000111;
        default: result = 8'b00000000;
    endcase
end

endmodule
